`define DIRECTION_READ	1'b0
`define DIRECTION_WRITE 1'b1

`define DIRECTION_READ	0x0
`define DIRECTION_WRITE 0x1
